`include "my_if.sv"
package my_exe_pkg;
    //`include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "my_driver.sv"
endpackage: my_exe_pkg
